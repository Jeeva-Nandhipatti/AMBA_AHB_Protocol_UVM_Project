//`include "uvm_macros.svh" 
package tb_pkg;
  `include "Seq_item.sv"
  `include "Sequence.sv"
  `include "Sequencer.sv"
  `include "Driver.sv"
  `include "Monitor.sv"
  `include "Agent.sv"
  `include "Scoreboard.sv"
  `include "Coverage.sv"
  `include "Environment.sv"
  `include "Test.sv"
endpackage
